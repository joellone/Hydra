module main;
    initial begin
        $display ("Hello iverilog");
        $finish;
    end
endmodule
